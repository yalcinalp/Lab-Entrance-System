`timescale 1ns / 1ps


module testbench;
	// Inputs
	reg I0;
	reg I1;
	reg I2;
	reg clk;
	// Outputs
	wire Q0;
	wire Q1;
	wire Z;

    // Result Memory
    reg[2:0] results0[7:0];
    reg[2:0] results1[7:0];
    reg[2:0] results2[7:0];
    // Scrambled Input Memory
    reg[2:0] scrInputs[7:0];
    reg[2:0] incInputs[7:0];
    reg[2:0] decInputs[7:0];
    // Loop iterator
    integer i;
    parameter INPUT_COMBINATIONS = 8;

	// Instantiate the Unit Under Test (UUT)
	ic1337 uut (.I0(I0),
                .I1(I1),
                .I2(I2),
                .clk(clk),
                .Q0(Q0),
                .Q1(Q1),
                .Z(Z));

    initial begin
        // Manually scramble inputs
        scrInputs[0] = 31'd2;
        scrInputs[1] = 31'd4;
        scrInputs[2] = 31'd6;
        scrInputs[3] = 31'd1;
        scrInputs[4] = 31'd0;
        scrInputs[5] = 31'd3;
        scrInputs[6] = 31'd7;
        scrInputs[7] = 31'd5;
        // Incrementing inputs
        incInputs[0] = 31'd0;
        incInputs[1] = 31'd1;
        incInputs[2] = 31'd2;
        incInputs[3] = 31'd3;
        incInputs[4] = 31'd4;
        incInputs[5] = 31'd5;
        incInputs[6] = 31'd6;
        incInputs[7] = 31'd7;
        // Decrementing inputs
        decInputs[0] = 31'd7;
        decInputs[1] = 31'd6;
        decInputs[2] = 31'd5;
        decInputs[3] = 31'd4;
        decInputs[4] = 31'd3;
        decInputs[5] = 31'd2;
        decInputs[6] = 31'd1;
        decInputs[7] = 31'd0;
        // Result list (generated by the code)
        results0[0] = 3'b000;
        results0[1] = 3'b000;
        results0[2] = 3'b000;
        results0[3] = 3'b110;
        results0[4] = 3'b011;
        results0[5] = 3'b011;
        results0[6] = 3'b011;
        results0[7] = 3'b011;
        //
        results1[0] = 3'b011;
        results1[1] = 3'b011;
        results1[2] = 3'b011;
        results1[3] = 3'b011;
        results1[4] = 3'b101;
        results1[5] = 3'b000;
        results1[6] = 3'b000;
        results1[7] = 3'b110;
        //
        results2[0] = 3'b000;
        results2[1] = 3'b011;
        results2[2] = 3'b011;
        results2[3] = 3'b101;
        results2[4] = 3'b011;
        results2[5] = 3'b101;
        results2[6] = 3'b101;
        results2[7] = 3'b101;
    end

    integer grade = 0;

    // Clock Related
    // At 5, 15, 25, .. clk will change 0->1
	// At 10, 20, 30, .. clk will change 1->0
    initial clk = 0;
    always #5 clk = ~clk;

	initial begin
        // (0ns) initialize I's just to be sure
        I0 = 1'b0;
        I1 = 1'b0;
        I2 = 1'b0;
        #6;
        // Enter to the loop after one ms later

        // Do a one round check of all bits
        // w/e it checks.

        //==========================//
        //         INCREMENT        //
        //==========================//
        // FOR LOOP SHOULD START 1NS AFTER POSEDGE CLOCK
        // Run the clock check the provided input with compared output
        for(i = 0; i < INPUT_COMBINATIONS; i = i + 1)
        begin
            // Time: (n + 1)
            // Decompose the i to bits
            I0 = incInputs[i][0];
            I1 = incInputs[i][1];
            I2 = incInputs[i][2];
            // Wait to next pos edge
            #10;
            $display("R = %b", {Z, Q1, Q0});
            // Check the output
            if(Q0 !== results0[i][0]) $display("Wrong Q0[%b], should be %b", Q0, results0[i][0]);
            else grade = grade + 1;
            if(Q1 !== results0[i][1]) $display("Wrong Q1[%b], should be %b", Q1, results0[i][1]);
            else grade = grade + 1;
            if( Z !== results0[i][2]) $display("Wrong  Z[%b], should be %b",  Z, results0[i][2]);
            else grade = grade + 1;
        end

        //==========================//
        //         DECREMENT        //
        //==========================//
        // FOR LOOP SHOULD START 1NS AFTER POSEDGE CLOCK
        // Run the clock check the provided input with compared output
        for(i = 0; i < INPUT_COMBINATIONS; i = i + 1)
        begin
            // Time: (n + 1)
            // Decompose the i to bits
            I0 = decInputs[i][0];
            I1 = decInputs[i][1];
            I2 = decInputs[i][2];
            // Wait to next pos edge
            #10;
            $display("R = %b", {Z, Q1, Q0});
            // Check the output
            if(Q0 !== results1[i][0]) $display("Wrong Q0[%b], should be %b", Q0, results1[i][0]);
            else grade = grade + 1;
            if(Q1 !== results1[i][1]) $display("Wrong Q1[%b], should be %b", Q1, results1[i][1]);
            else grade = grade + 1;
            if( Z !== results1[i][2]) $display("Wrong  Z[%b], should be %b",  Z, results1[i][2]);
            else grade = grade + 1;
        end

        //==========================//
        //         SCRAMBLED        //
        //==========================//
        // FOR LOOP SHOULD START 1NS AFTER POSEDGE CLOCK
        // Run the clock check the provided input with compared output
        for(i = 0; i < INPUT_COMBINATIONS; i = i + 1)
        begin
            // Time: (n + 1)
            // Decompose the i to bits
            I0 = scrInputs[i][0];
            I1 = scrInputs[i][1];
            I2 = scrInputs[i][2];
            // Wait to next pos edge
            #10;
            $display("R = %b", {Z, Q1, Q0});
            // Check the output
            if(Q0 !== results2[i][0]) $display("Wrong Q0[%b], should be %b", Q0, results2[i][0]);
            else grade = grade + 1;
            if(Q1 !== results2[i][1]) $display("Wrong Q1[%b], should be %b", Q1, results2[i][1]);
            else grade = grade + 1;
            if( Z !== results2[i][2]) $display("Wrong  Z[%b], should be %b",  Z, results2[i][2]);
            else grade = grade + 1;
        end
        #1
        $display("Result is:%d", grade);
		$finish;
	end

endmodule

